-------------------------------------------------------------------------------
--
-- Title       : alu
-- Design      : test
-- Author      : test
-- Company     : Test
--
-------------------------------------------------------------------------------
--
-- File        : C:\My_Designs\architecturelab\test\src\alu.vhd
-- Generated   : Wed Dec 11 14:43:25 2024
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {alu} architecture {alu}}



entity alu is
end alu;

--}} End of automatically maintained section

architecture alu of alu is
begin

	 -- enter your statements here --

end alu;
